module vitrine

// TODO: This needn't be public
pub struct Resolved {
  pub mut:
    size Vector2
    position Vector2
}