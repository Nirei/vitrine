module vitrine

struct Resolved {
pub mut:
	size     Vector2
	position Vector2
}
